// -----------------------------------------------------------------------------
// GHASH subkey generator: computes H = AES(K, 0^128) whenever a new key arrives
// Supports optional sharing of an external aes_core instance.
// -----------------------------------------------------------------------------
module h_subkey #(
    parameter SHARED_AES = 0
) (
    input  wire         clk,
    input  wire         rst_n,
    input  wire [255:0] key_in,
    input  wire         key_we,
    input  wire         aes256_en,
    output wire [127:0] H,
    output wire         H_valid,
    // Shared AES interface (used when SHARED_AES != 0)
    output wire         aes_req,
    input  wire         aes_gnt,
    output wire         aes_init,
    output wire         aes_next,
    output wire [255:0] aes_key,
    output wire         aes_keylen,
    output wire [127:0] aes_block,
    input  wire         aes_ready,
    input  wire [127:0] aes_result,
    input  wire         aes_result_valid
);

    localparam ST_IDLE       = 3'd0;
    localparam ST_ISSUE_INIT = 3'd1;
    localparam ST_WAIT_INIT  = 3'd2;
    localparam ST_ISSUE_NEXT = 3'd3;
    localparam ST_WAIT_RES   = 3'd4;

    reg [2:0]   state_reg;
    reg [2:0]   state_next;

    reg [255:0] key_active_reg;
    reg [255:0] key_active_next;
    reg         keylen_active_reg;
    reg         keylen_active_next;

    reg [255:0] key_queue_reg;
    reg [255:0] key_queue_next;
    reg         keylen_queue_reg;
    reg         keylen_queue_next;
    reg         queue_valid_reg;
    reg         queue_valid_next;

    reg         compute_pending_reg;
    reg         compute_pending_next;

    reg [127:0] h_reg;
    reg [127:0] h_next;
    reg         h_valid_reg;
    reg         h_valid_next;

    wire [255:0] sanitized_key    = aes256_en ? key_in : {128'h0, key_in[127:0]};
    wire         sanitized_keylen = aes256_en;

    wire         have_grant = (SHARED_AES != 0) ? aes_gnt : 1'b1;

    wire         core_init = (state_reg == ST_ISSUE_INIT);
    wire         core_next = (state_reg == ST_ISSUE_NEXT);

    wire         core_ready;
    wire [127:0] core_result;
    wire         core_result_valid;

    assign H       = h_reg;
    assign H_valid = h_valid_reg;

    assign aes_block = 128'h0;
    assign aes_key   = (SHARED_AES != 0) ? key_active_reg : 256'h0;
    assign aes_keylen = (SHARED_AES != 0) ? keylen_active_reg : 1'b0;
    assign aes_init  = (SHARED_AES != 0) ? core_init : 1'b0;
    assign aes_next  = (SHARED_AES != 0) ? core_next : 1'b0;
    assign aes_req   = (SHARED_AES != 0) ? (queue_valid_reg | compute_pending_reg | (state_reg != ST_IDLE)) : 1'b0;

    // ------------------------------------------------------------------
    // Sequential registers
    // ------------------------------------------------------------------
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state_reg            <= ST_IDLE;
            key_active_reg       <= 256'h0;
            keylen_active_reg    <= 1'b0;
            key_queue_reg        <= 256'h0;
            keylen_queue_reg     <= 1'b0;
            queue_valid_reg      <= 1'b0;
            compute_pending_reg  <= 1'b0;
            h_reg                <= 128'h0;
            h_valid_reg          <= 1'b0;
        end else begin
            state_reg            <= state_next;
            key_active_reg       <= key_active_next;
            keylen_active_reg    <= keylen_active_next;
            key_queue_reg        <= key_queue_next;
            keylen_queue_reg     <= keylen_queue_next;
            queue_valid_reg      <= queue_valid_next;
            compute_pending_reg  <= compute_pending_next;
            h_reg                <= h_next;
            h_valid_reg          <= h_valid_next;
        end
    end

    // ------------------------------------------------------------------
    // Combinational control
    // ------------------------------------------------------------------
    always @* begin
        state_next            = state_reg;
        key_active_next       = key_active_reg;
        keylen_active_next    = keylen_active_reg;
        key_queue_next        = key_queue_reg;
        keylen_queue_next     = keylen_queue_reg;
        queue_valid_next      = queue_valid_reg;
        compute_pending_next  = compute_pending_reg;
        h_next                = h_reg;
        h_valid_next          = 1'b0;

        // Promote queued key when idle and no pending compute
        if ((state_reg == ST_IDLE) && !compute_pending_next && queue_valid_reg) begin
            key_active_next      = key_queue_reg;
            keylen_active_next   = keylen_queue_reg;
            compute_pending_next = 1'b1;
            queue_valid_next     = 1'b0;
        end

        // Capture new key writes
        if (key_we) begin
            if ((state_reg == ST_IDLE) && !compute_pending_next) begin
                key_active_next      = sanitized_key;
                keylen_active_next   = sanitized_keylen;
                compute_pending_next = 1'b1;
            end else begin
                key_queue_next    = sanitized_key;
                keylen_queue_next = sanitized_keylen;
                queue_valid_next  = 1'b1;
            end
        end

        case (state_reg)
            ST_IDLE: begin
                if (compute_pending_next && have_grant) begin
                    state_next           = ST_ISSUE_INIT;
                    compute_pending_next = 1'b0;
                end
            end

            ST_ISSUE_INIT: begin
                state_next = ST_WAIT_INIT;
            end

            ST_WAIT_INIT: begin
                if (core_ready) begin
                    state_next = ST_ISSUE_NEXT;
                end
            end

            ST_ISSUE_NEXT: begin
                state_next = ST_WAIT_RES;
            end

            ST_WAIT_RES: begin
                if (core_result_valid) begin
                    h_next       = core_result;
                    h_valid_next = 1'b1;

                    if (queue_valid_reg) begin
                        key_active_next      = key_queue_reg;
                        keylen_active_next   = keylen_queue_reg;
                        queue_valid_next     = 1'b0;
                        compute_pending_next = 1'b1;
                    end

                    state_next = ST_IDLE;
                end
            end

            default: begin
                state_next = ST_IDLE;
            end
        endcase
    end

    // ------------------------------------------------------------------
    // AES core hookup (internal or shared)
    // ------------------------------------------------------------------
    wire        core_ready_int;
    wire [127:0] core_result_int;
    wire        core_result_valid_int;

    generate
        if (SHARED_AES == 0) begin : gen_internal_aes
            aes_core u_aes_core (
                .clk          (clk),
                .reset_n      (rst_n),
                .encdec       (1'b1),
                .init         (core_init),
                .next         (core_next),
                .ready        (core_ready_int),
                .key          (key_active_reg),
                .keylen       (keylen_active_reg),
                .block        (128'h0),
                .result       (core_result_int),
                .result_valid (core_result_valid_int)
            );
        end else begin : gen_shared_aes
            assign core_ready_int        = 1'b0;
            assign core_result_int       = 128'h0;
            assign core_result_valid_int = 1'b0;
        end
    endgenerate

    assign core_ready        = (SHARED_AES == 0) ? core_ready_int : aes_ready;
    assign core_result       = (SHARED_AES == 0) ? core_result_int : aes_result;
    assign core_result_valid = (SHARED_AES == 0) ? core_result_valid_int : aes_result_valid;

endmodule



